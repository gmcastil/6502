module alu
  #(
    // parameter
    )
   (
    input A,
    input B,
    input carry_in,
    output overflow,
    output carry,
    output half_carry
